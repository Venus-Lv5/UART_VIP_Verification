`ifndef GUARD_UART_TEST_PKG__SV
`define GUARD_UART_TEST_PKG__SV


package test_pkg;
	import uvm_pkg::*;
	import ahb_pkg::*;
	import env_pkg::*;
	import seq_pkg::*;
	import uart_regmodel_pkg::*;
	import uart_pkg::*;

	`include "uart_base_test.sv"

	`include "reg_rsvd_test.sv"
	`include "reg_rw_test.sv"
	`include "reg_default_test.sv"
	`include "reg_w1c_test.sv"
	
	`include "x13_2400_test.sv"
	`include "x13_4800_test.sv"
	`include "x13_9600_test.sv"
	`include "x13_19200_test.sv"
	`include "x13_38400_test.sv"
	`include "x13_76800_test.sv"
	`include "x13_115200_test.sv"
	`include "x13_custom_test.sv"

	`include "x16_2400_test.sv"
	`include "x16_4800_test.sv"
	`include "x16_9600_test.sv"
	`include "x16_19200_test.sv"
	`include "x16_38400_test.sv"
	`include "x16_76800_test.sv"
	`include "x16_115200_test.sv"
	`include "x16_custom_test.sv"

	`include "transmit_2400_5_none_1_test.sv"
	`include "transmit_2400_5_none_2_test.sv"
	`include "transmit_2400_5_odd_1_test.sv"
	`include "transmit_2400_5_odd_2_test.sv"
	`include "transmit_2400_5_even_1_test.sv"
	`include "transmit_2400_5_even_2_test.sv"

	`include "transmit_2400_6_none_1_test.sv"
	`include "transmit_2400_6_none_2_test.sv"
	`include "transmit_2400_6_odd_1_test.sv"
	`include "transmit_2400_6_odd_2_test.sv"
	`include "transmit_2400_6_even_1_test.sv"
	`include "transmit_2400_6_even_2_test.sv"
	
	`include "transmit_2400_7_none_1_test.sv"
	`include "transmit_2400_7_none_2_test.sv"
	`include "transmit_2400_7_odd_1_test.sv"
	`include "transmit_2400_7_odd_2_test.sv"
	`include "transmit_2400_7_even_1_test.sv"
	`include "transmit_2400_7_even_2_test.sv"
	
	`include "transmit_2400_8_none_1_test.sv"
	`include "transmit_2400_8_none_2_test.sv"
	`include "transmit_2400_8_odd_1_test.sv"
	`include "transmit_2400_8_odd_2_test.sv"
	`include "transmit_2400_8_even_1_test.sv"
	`include "transmit_2400_8_even_2_test.sv"
	
	`include "transmit_4800_5_none_1_test.sv"
	`include "transmit_4800_5_none_2_test.sv"
	`include "transmit_4800_5_odd_1_test.sv"
	`include "transmit_4800_5_odd_2_test.sv"
	`include "transmit_4800_5_even_1_test.sv"
	`include "transmit_4800_5_even_2_test.sv"

	`include "transmit_4800_6_none_1_test.sv"
	`include "transmit_4800_6_none_2_test.sv"
	`include "transmit_4800_6_odd_1_test.sv"
	`include "transmit_4800_6_odd_2_test.sv"
	`include "transmit_4800_6_even_1_test.sv"
	`include "transmit_4800_6_even_2_test.sv"
	
	`include "transmit_4800_7_none_1_test.sv"
	`include "transmit_4800_7_none_2_test.sv"
	`include "transmit_4800_7_odd_1_test.sv"
	`include "transmit_4800_7_odd_2_test.sv"
	`include "transmit_4800_7_even_1_test.sv"
	`include "transmit_4800_7_even_2_test.sv"
	
	`include "transmit_4800_8_none_1_test.sv"
	`include "transmit_4800_8_none_2_test.sv"
	`include "transmit_4800_8_odd_1_test.sv"
	`include "transmit_4800_8_odd_2_test.sv"
	`include "transmit_4800_8_even_1_test.sv"
	`include "transmit_4800_8_even_2_test.sv"
	
	`include "transmit_9600_5_none_1_test.sv"
	`include "transmit_9600_5_none_2_test.sv"
	`include "transmit_9600_5_odd_1_test.sv"
	`include "transmit_9600_5_odd_2_test.sv"
	`include "transmit_9600_5_even_1_test.sv"
	`include "transmit_9600_5_even_2_test.sv"

	`include "transmit_9600_6_none_1_test.sv"
	`include "transmit_9600_6_none_2_test.sv"
	`include "transmit_9600_6_odd_1_test.sv"
	`include "transmit_9600_6_odd_2_test.sv"
	`include "transmit_9600_6_even_1_test.sv"
	`include "transmit_9600_6_even_2_test.sv"
	
	`include "transmit_9600_7_none_1_test.sv"
	`include "transmit_9600_7_none_2_test.sv"
	`include "transmit_9600_7_odd_1_test.sv"
	`include "transmit_9600_7_odd_2_test.sv"
	`include "transmit_9600_7_even_1_test.sv"
	`include "transmit_9600_7_even_2_test.sv"
	
	`include "transmit_9600_8_none_1_test.sv"
	`include "transmit_9600_8_none_2_test.sv"
	`include "transmit_9600_8_odd_1_test.sv"
	`include "transmit_9600_8_odd_2_test.sv"
	`include "transmit_9600_8_even_1_test.sv"
	`include "transmit_9600_8_even_2_test.sv"
	
	`include "transmit_19200_5_none_1_test.sv"
	`include "transmit_19200_5_none_2_test.sv"
	`include "transmit_19200_5_odd_1_test.sv"
	`include "transmit_19200_5_odd_2_test.sv"
	`include "transmit_19200_5_even_1_test.sv"
	`include "transmit_19200_5_even_2_test.sv"

	`include "transmit_19200_6_none_1_test.sv"
	`include "transmit_19200_6_none_2_test.sv"
	`include "transmit_19200_6_odd_1_test.sv"
	`include "transmit_19200_6_odd_2_test.sv"
	`include "transmit_19200_6_even_1_test.sv"
	`include "transmit_19200_6_even_2_test.sv"
	
	`include "transmit_19200_7_none_1_test.sv"
	`include "transmit_19200_7_none_2_test.sv"
	`include "transmit_19200_7_odd_1_test.sv"
	`include "transmit_19200_7_odd_2_test.sv"
	`include "transmit_19200_7_even_1_test.sv"
	`include "transmit_19200_7_even_2_test.sv"
	
	`include "transmit_19200_8_none_1_test.sv"
	`include "transmit_19200_8_none_2_test.sv"
	`include "transmit_19200_8_odd_1_test.sv"
	`include "transmit_19200_8_odd_2_test.sv"
	`include "transmit_19200_8_even_1_test.sv"
	`include "transmit_19200_8_even_2_test.sv"
	
	`include "transmit_38400_5_none_1_test.sv"
	`include "transmit_38400_5_none_2_test.sv"
	`include "transmit_38400_5_odd_1_test.sv"
	`include "transmit_38400_5_odd_2_test.sv"
	`include "transmit_38400_5_even_1_test.sv"
	`include "transmit_38400_5_even_2_test.sv"

	`include "transmit_38400_6_none_1_test.sv"
	`include "transmit_38400_6_none_2_test.sv"
	`include "transmit_38400_6_odd_1_test.sv"
	`include "transmit_38400_6_odd_2_test.sv"
	`include "transmit_38400_6_even_1_test.sv"
	`include "transmit_38400_6_even_2_test.sv"
	
	`include "transmit_38400_7_none_1_test.sv"
	`include "transmit_38400_7_none_2_test.sv"
	`include "transmit_38400_7_odd_1_test.sv"
	`include "transmit_38400_7_odd_2_test.sv"
	`include "transmit_38400_7_even_1_test.sv"
	`include "transmit_38400_7_even_2_test.sv"
	
	`include "transmit_38400_8_none_1_test.sv"
	`include "transmit_38400_8_none_2_test.sv"
	`include "transmit_38400_8_odd_1_test.sv"
	`include "transmit_38400_8_odd_2_test.sv"
	`include "transmit_38400_8_even_1_test.sv"
	`include "transmit_38400_8_even_2_test.sv"
	
	`include "transmit_76800_5_none_1_test.sv"
	`include "transmit_76800_5_none_2_test.sv"
	`include "transmit_76800_5_odd_1_test.sv"
	`include "transmit_76800_5_odd_2_test.sv"
	`include "transmit_76800_5_even_1_test.sv"
	`include "transmit_76800_5_even_2_test.sv"

	`include "transmit_76800_6_none_1_test.sv"
	`include "transmit_76800_6_none_2_test.sv"
	`include "transmit_76800_6_odd_1_test.sv"
	`include "transmit_76800_6_odd_2_test.sv"
	`include "transmit_76800_6_even_1_test.sv"
	`include "transmit_76800_6_even_2_test.sv"
	
	`include "transmit_76800_7_none_1_test.sv"
	`include "transmit_76800_7_none_2_test.sv"
	`include "transmit_76800_7_odd_1_test.sv"
	`include "transmit_76800_7_odd_2_test.sv"
	`include "transmit_76800_7_even_1_test.sv"
	`include "transmit_76800_7_even_2_test.sv"
	
	`include "transmit_76800_8_none_1_test.sv"
	`include "transmit_76800_8_none_2_test.sv"
	`include "transmit_76800_8_odd_1_test.sv"
	`include "transmit_76800_8_odd_2_test.sv"
	`include "transmit_76800_8_even_1_test.sv"
	`include "transmit_76800_8_even_2_test.sv"
	
	`include "transmit_115200_5_none_1_test.sv"
	`include "transmit_115200_5_none_2_test.sv"
	`include "transmit_115200_5_odd_1_test.sv"
	`include "transmit_115200_5_odd_2_test.sv"
	`include "transmit_115200_5_even_1_test.sv"
	`include "transmit_115200_5_even_2_test.sv"

	`include "transmit_115200_6_none_1_test.sv"
	`include "transmit_115200_6_none_2_test.sv"
	`include "transmit_115200_6_odd_1_test.sv"
	`include "transmit_115200_6_odd_2_test.sv"
	`include "transmit_115200_6_even_1_test.sv"
	`include "transmit_115200_6_even_2_test.sv"
	
	`include "transmit_115200_7_none_1_test.sv"
	`include "transmit_115200_7_none_2_test.sv"
	`include "transmit_115200_7_odd_1_test.sv"
	`include "transmit_115200_7_odd_2_test.sv"
	`include "transmit_115200_7_even_1_test.sv"
	`include "transmit_115200_7_even_2_test.sv"
	
	`include "transmit_115200_8_none_1_test.sv"
	`include "transmit_115200_8_none_2_test.sv"
	`include "transmit_115200_8_odd_1_test.sv"
	`include "transmit_115200_8_odd_2_test.sv"
	`include "transmit_115200_8_even_1_test.sv"
	`include "transmit_115200_8_even_2_test.sv"
	
	`include "transmit_custom_5_none_1_test.sv"
	`include "transmit_custom_5_none_2_test.sv"
	`include "transmit_custom_5_odd_1_test.sv"
	`include "transmit_custom_5_odd_2_test.sv"
	`include "transmit_custom_5_even_1_test.sv"
	`include "transmit_custom_5_even_2_test.sv"

	`include "transmit_custom_6_none_1_test.sv"
	`include "transmit_custom_6_none_2_test.sv"
	`include "transmit_custom_6_odd_1_test.sv"
	`include "transmit_custom_6_odd_2_test.sv"
	`include "transmit_custom_6_even_1_test.sv"
	`include "transmit_custom_6_even_2_test.sv"
	
	`include "transmit_custom_7_none_1_test.sv"
	`include "transmit_custom_7_none_2_test.sv"
	`include "transmit_custom_7_odd_1_test.sv"
	`include "transmit_custom_7_odd_2_test.sv"
	`include "transmit_custom_7_even_1_test.sv"
	`include "transmit_custom_7_even_2_test.sv"
	
	`include "transmit_custom_8_none_1_test.sv"
	`include "transmit_custom_8_none_2_test.sv"
	`include "transmit_custom_8_odd_1_test.sv"
	`include "transmit_custom_8_odd_2_test.sv"
	`include "transmit_custom_8_even_1_test.sv"
	`include "transmit_custom_8_even_2_test.sv"

	`include "transmit_dynamic_config_test.sv"



	`include "receive_2400_5_none_1_test.sv"
	`include "receive_2400_5_none_2_test.sv"
	`include "receive_2400_5_odd_1_test.sv"
	`include "receive_2400_5_odd_2_test.sv"
	`include "receive_2400_5_even_1_test.sv"
	`include "receive_2400_5_even_2_test.sv"

	`include "receive_2400_6_none_1_test.sv"
	`include "receive_2400_6_none_2_test.sv"
	`include "receive_2400_6_odd_1_test.sv"
	`include "receive_2400_6_odd_2_test.sv"
	`include "receive_2400_6_even_1_test.sv"
	`include "receive_2400_6_even_2_test.sv"

	`include "receive_2400_7_none_1_test.sv"
	`include "receive_2400_7_none_2_test.sv"
	`include "receive_2400_7_odd_1_test.sv"
	`include "receive_2400_7_odd_2_test.sv"
	`include "receive_2400_7_even_1_test.sv"
	`include "receive_2400_7_even_2_test.sv"

	`include "receive_2400_8_none_1_test.sv"
	`include "receive_2400_8_none_2_test.sv"
	`include "receive_2400_8_odd_1_test.sv"
	`include "receive_2400_8_odd_2_test.sv"
	`include "receive_2400_8_even_1_test.sv"
	`include "receive_2400_8_even_2_test.sv"

	`include "receive_4800_5_none_1_test.sv"
	`include "receive_4800_5_none_2_test.sv"
	`include "receive_4800_5_odd_1_test.sv"
	`include "receive_4800_5_odd_2_test.sv"
	`include "receive_4800_5_even_1_test.sv"
	`include "receive_4800_5_even_2_test.sv"

	`include "receive_4800_6_none_1_test.sv"
	`include "receive_4800_6_none_2_test.sv"
	`include "receive_4800_6_odd_1_test.sv"
	`include "receive_4800_6_odd_2_test.sv"
	`include "receive_4800_6_even_1_test.sv"
	`include "receive_4800_6_even_2_test.sv"

	`include "receive_4800_7_none_1_test.sv"
	`include "receive_4800_7_none_2_test.sv"
	`include "receive_4800_7_odd_1_test.sv"
	`include "receive_4800_7_odd_2_test.sv"
	`include "receive_4800_7_even_1_test.sv"
	`include "receive_4800_7_even_2_test.sv"

	`include "receive_4800_8_none_1_test.sv"
	`include "receive_4800_8_none_2_test.sv"
	`include "receive_4800_8_odd_1_test.sv"
	`include "receive_4800_8_odd_2_test.sv"
	`include "receive_4800_8_even_1_test.sv"
	`include "receive_4800_8_even_2_test.sv"

	`include "receive_9600_5_none_1_test.sv"
	`include "receive_9600_5_none_2_test.sv"
	`include "receive_9600_5_odd_1_test.sv"
	`include "receive_9600_5_odd_2_test.sv"
	`include "receive_9600_5_even_1_test.sv"
	`include "receive_9600_5_even_2_test.sv"

	`include "receive_9600_6_none_1_test.sv"
	`include "receive_9600_6_none_2_test.sv"
	`include "receive_9600_6_odd_1_test.sv"
	`include "receive_9600_6_odd_2_test.sv"
	`include "receive_9600_6_even_1_test.sv"
	`include "receive_9600_6_even_2_test.sv"

	`include "receive_9600_7_none_1_test.sv"
	`include "receive_9600_7_none_2_test.sv"
	`include "receive_9600_7_odd_1_test.sv"
	`include "receive_9600_7_odd_2_test.sv"
	`include "receive_9600_7_even_1_test.sv"
	`include "receive_9600_7_even_2_test.sv"

	`include "receive_9600_8_none_1_test.sv"
	`include "receive_9600_8_none_2_test.sv"
	`include "receive_9600_8_odd_1_test.sv"
	`include "receive_9600_8_odd_2_test.sv"
	`include "receive_9600_8_even_1_test.sv"
	`include "receive_9600_8_even_2_test.sv"

	`include "receive_19200_5_none_1_test.sv"
	`include "receive_19200_5_none_2_test.sv"
	`include "receive_19200_5_odd_1_test.sv"
	`include "receive_19200_5_odd_2_test.sv"
	`include "receive_19200_5_even_1_test.sv"
	`include "receive_19200_5_even_2_test.sv"

	`include "receive_19200_6_none_1_test.sv"
	`include "receive_19200_6_none_2_test.sv"
	`include "receive_19200_6_odd_1_test.sv"
	`include "receive_19200_6_odd_2_test.sv"
	`include "receive_19200_6_even_1_test.sv"
	`include "receive_19200_6_even_2_test.sv"

	`include "receive_19200_7_none_1_test.sv"
	`include "receive_19200_7_none_2_test.sv"
	`include "receive_19200_7_odd_1_test.sv"
	`include "receive_19200_7_odd_2_test.sv"
	`include "receive_19200_7_even_1_test.sv"
	`include "receive_19200_7_even_2_test.sv"

	`include "receive_19200_8_none_1_test.sv"
	`include "receive_19200_8_none_2_test.sv"
	`include "receive_19200_8_odd_1_test.sv"
	`include "receive_19200_8_odd_2_test.sv"
	`include "receive_19200_8_even_1_test.sv"
	`include "receive_19200_8_even_2_test.sv"

	`include "receive_38400_5_none_1_test.sv"
	`include "receive_38400_5_none_2_test.sv"
	`include "receive_38400_5_odd_1_test.sv"
	`include "receive_38400_5_odd_2_test.sv"
	`include "receive_38400_5_even_1_test.sv"
	`include "receive_38400_5_even_2_test.sv"

	`include "receive_38400_6_none_1_test.sv"
	`include "receive_38400_6_none_2_test.sv"
	`include "receive_38400_6_odd_1_test.sv"
	`include "receive_38400_6_odd_2_test.sv"
	`include "receive_38400_6_even_1_test.sv"
	`include "receive_38400_6_even_2_test.sv"

	`include "receive_38400_7_none_1_test.sv"
	`include "receive_38400_7_none_2_test.sv"
	`include "receive_38400_7_odd_1_test.sv"
	`include "receive_38400_7_odd_2_test.sv"
	`include "receive_38400_7_even_1_test.sv"
	`include "receive_38400_7_even_2_test.sv"

	`include "receive_38400_8_none_1_test.sv"
	`include "receive_38400_8_none_2_test.sv"
	`include "receive_38400_8_odd_1_test.sv"
	`include "receive_38400_8_odd_2_test.sv"
	`include "receive_38400_8_even_1_test.sv"
	`include "receive_38400_8_even_2_test.sv"

	`include "receive_76800_5_none_1_test.sv"
	`include "receive_76800_5_none_2_test.sv"
	`include "receive_76800_5_odd_1_test.sv"
	`include "receive_76800_5_odd_2_test.sv"
	`include "receive_76800_5_even_1_test.sv"
	`include "receive_76800_5_even_2_test.sv"

	`include "receive_76800_6_none_1_test.sv"
	`include "receive_76800_6_none_2_test.sv"
	`include "receive_76800_6_odd_1_test.sv"
	`include "receive_76800_6_odd_2_test.sv"
	`include "receive_76800_6_even_1_test.sv"
	`include "receive_76800_6_even_2_test.sv"

	`include "receive_76800_7_none_1_test.sv"
	`include "receive_76800_7_none_2_test.sv"
	`include "receive_76800_7_odd_1_test.sv"
	`include "receive_76800_7_odd_2_test.sv"
	`include "receive_76800_7_even_1_test.sv"
	`include "receive_76800_7_even_2_test.sv"

	`include "receive_76800_8_none_1_test.sv"
	`include "receive_76800_8_none_2_test.sv"
	`include "receive_76800_8_odd_1_test.sv"
	`include "receive_76800_8_odd_2_test.sv"
	`include "receive_76800_8_even_1_test.sv"
	`include "receive_76800_8_even_2_test.sv"

	`include "receive_115200_5_none_1_test.sv"
	`include "receive_115200_5_none_2_test.sv"
	`include "receive_115200_5_odd_1_test.sv"
	`include "receive_115200_5_odd_2_test.sv"
	`include "receive_115200_5_even_1_test.sv"
	`include "receive_115200_5_even_2_test.sv"

	`include "receive_115200_6_none_1_test.sv"
	`include "receive_115200_6_none_2_test.sv"
	`include "receive_115200_6_odd_1_test.sv"
	`include "receive_115200_6_odd_2_test.sv"
	`include "receive_115200_6_even_1_test.sv"
	`include "receive_115200_6_even_2_test.sv"

	`include "receive_115200_7_none_1_test.sv"
	`include "receive_115200_7_none_2_test.sv"
	`include "receive_115200_7_odd_1_test.sv"
	`include "receive_115200_7_odd_2_test.sv"
	`include "receive_115200_7_even_1_test.sv"
	`include "receive_115200_7_even_2_test.sv"

	`include "receive_115200_8_none_1_test.sv"
	`include "receive_115200_8_none_2_test.sv"
	`include "receive_115200_8_odd_1_test.sv"
	`include "receive_115200_8_odd_2_test.sv"
	`include "receive_115200_8_even_1_test.sv"
	`include "receive_115200_8_even_2_test.sv"

	`include "receive_custom_5_none_1_test.sv"
	`include "receive_custom_5_none_2_test.sv"
	`include "receive_custom_5_odd_1_test.sv"
	`include "receive_custom_5_odd_2_test.sv"
	`include "receive_custom_5_even_1_test.sv"
	`include "receive_custom_5_even_2_test.sv"

	`include "receive_custom_6_none_1_test.sv"
	`include "receive_custom_6_none_2_test.sv"
	`include "receive_custom_6_odd_1_test.sv"
	`include "receive_custom_6_odd_2_test.sv"
	`include "receive_custom_6_even_1_test.sv"
	`include "receive_custom_6_even_2_test.sv"

	`include "receive_custom_7_none_1_test.sv"
	`include "receive_custom_7_none_2_test.sv"
	`include "receive_custom_7_odd_1_test.sv"
	`include "receive_custom_7_odd_2_test.sv"
	`include "receive_custom_7_even_1_test.sv"
	`include "receive_custom_7_even_2_test.sv"

	`include "receive_custom_8_none_1_test.sv"
	`include "receive_custom_8_none_2_test.sv"
	`include "receive_custom_8_odd_1_test.sv"
	`include "receive_custom_8_odd_2_test.sv"
	`include "receive_custom_8_even_1_test.sv"
	`include "receive_custom_8_even_2_test.sv"

	`include "receive_dynamic_config_test.sv"

	`include "full_2400_5_none_1_test.sv"
	`include "full_2400_5_none_2_test.sv"
	`include "full_2400_5_odd_1_test.sv"
	`include "full_2400_5_odd_2_test.sv"
	`include "full_2400_5_even_1_test.sv"
	`include "full_2400_5_even_2_test.sv"

	`include "full_2400_6_none_1_test.sv"
	`include "full_2400_6_none_2_test.sv"
	`include "full_2400_6_odd_1_test.sv"
	`include "full_2400_6_odd_2_test.sv"
	`include "full_2400_6_even_1_test.sv"
	`include "full_2400_6_even_2_test.sv"

	`include "full_2400_7_none_1_test.sv"
	`include "full_2400_7_none_2_test.sv"
	`include "full_2400_7_odd_1_test.sv"
	`include "full_2400_7_odd_2_test.sv"
	`include "full_2400_7_even_1_test.sv"
	`include "full_2400_7_even_2_test.sv"

	`include "full_2400_8_none_1_test.sv"
	`include "full_2400_8_none_2_test.sv"
	`include "full_2400_8_odd_1_test.sv"
	`include "full_2400_8_odd_2_test.sv"
	`include "full_2400_8_even_1_test.sv"
	`include "full_2400_8_even_2_test.sv"

	`include "full_4800_5_none_1_test.sv"
	`include "full_4800_5_none_2_test.sv"
	`include "full_4800_5_odd_1_test.sv"
	`include "full_4800_5_odd_2_test.sv"
	`include "full_4800_5_even_1_test.sv"
	`include "full_4800_5_even_2_test.sv"

	`include "full_4800_6_none_1_test.sv"
	`include "full_4800_6_none_2_test.sv"
	`include "full_4800_6_odd_1_test.sv"
	`include "full_4800_6_odd_2_test.sv"
	`include "full_4800_6_even_1_test.sv"
	`include "full_4800_6_even_2_test.sv"

	`include "full_4800_7_none_1_test.sv"
	`include "full_4800_7_none_2_test.sv"
	`include "full_4800_7_odd_1_test.sv"
	`include "full_4800_7_odd_2_test.sv"
	`include "full_4800_7_even_1_test.sv"
	`include "full_4800_7_even_2_test.sv"

	`include "full_4800_8_none_1_test.sv"
	`include "full_4800_8_none_2_test.sv"
	`include "full_4800_8_odd_1_test.sv"
	`include "full_4800_8_odd_2_test.sv"
	`include "full_4800_8_even_1_test.sv"
	`include "full_4800_8_even_2_test.sv"

	`include "full_9600_5_none_1_test.sv"
	`include "full_9600_5_none_2_test.sv"
	`include "full_9600_5_odd_1_test.sv"
	`include "full_9600_5_odd_2_test.sv"
	`include "full_9600_5_even_1_test.sv"
	`include "full_9600_5_even_2_test.sv"

	`include "full_9600_6_none_1_test.sv"
	`include "full_9600_6_none_2_test.sv"
	`include "full_9600_6_odd_1_test.sv"
	`include "full_9600_6_odd_2_test.sv"
	`include "full_9600_6_even_1_test.sv"
	`include "full_9600_6_even_2_test.sv"

	`include "full_9600_7_none_1_test.sv"
	`include "full_9600_7_none_2_test.sv"
	`include "full_9600_7_odd_1_test.sv"
	`include "full_9600_7_odd_2_test.sv"
	`include "full_9600_7_even_1_test.sv"
	`include "full_9600_7_even_2_test.sv"

	`include "full_9600_8_none_1_test.sv"
	`include "full_9600_8_none_2_test.sv"
	`include "full_9600_8_odd_1_test.sv"
	`include "full_9600_8_odd_2_test.sv"
	`include "full_9600_8_even_1_test.sv"
	`include "full_9600_8_even_2_test.sv"

	`include "full_19200_5_none_1_test.sv"
	`include "full_19200_5_none_2_test.sv"
	`include "full_19200_5_odd_1_test.sv"
	`include "full_19200_5_odd_2_test.sv"
	`include "full_19200_5_even_1_test.sv"
	`include "full_19200_5_even_2_test.sv"

	`include "full_19200_6_none_1_test.sv"
	`include "full_19200_6_none_2_test.sv"
	`include "full_19200_6_odd_1_test.sv"
	`include "full_19200_6_odd_2_test.sv"
	`include "full_19200_6_even_1_test.sv"
	`include "full_19200_6_even_2_test.sv"

	`include "full_19200_7_none_1_test.sv"
	`include "full_19200_7_none_2_test.sv"
	`include "full_19200_7_odd_1_test.sv"
	`include "full_19200_7_odd_2_test.sv"
	`include "full_19200_7_even_1_test.sv"
	`include "full_19200_7_even_2_test.sv"

	`include "full_19200_8_none_1_test.sv"
	`include "full_19200_8_none_2_test.sv"
	`include "full_19200_8_odd_1_test.sv"
	`include "full_19200_8_odd_2_test.sv"
	`include "full_19200_8_even_1_test.sv"
	`include "full_19200_8_even_2_test.sv"

	`include "full_38400_5_none_1_test.sv"
	`include "full_38400_5_none_2_test.sv"
	`include "full_38400_5_odd_1_test.sv"
	`include "full_38400_5_odd_2_test.sv"
	`include "full_38400_5_even_1_test.sv"
	`include "full_38400_5_even_2_test.sv"

	`include "full_38400_6_none_1_test.sv"
	`include "full_38400_6_none_2_test.sv"
	`include "full_38400_6_odd_1_test.sv"
	`include "full_38400_6_odd_2_test.sv"
	`include "full_38400_6_even_1_test.sv"
	`include "full_38400_6_even_2_test.sv"

	`include "full_38400_7_none_1_test.sv"
	`include "full_38400_7_none_2_test.sv"
	`include "full_38400_7_odd_1_test.sv"
	`include "full_38400_7_odd_2_test.sv"
	`include "full_38400_7_even_1_test.sv"
	`include "full_38400_7_even_2_test.sv"

	`include "full_38400_8_none_1_test.sv"
	`include "full_38400_8_none_2_test.sv"
	`include "full_38400_8_odd_1_test.sv"
	`include "full_38400_8_odd_2_test.sv"
	`include "full_38400_8_even_1_test.sv"
	`include "full_38400_8_even_2_test.sv"

	`include "full_76800_5_none_1_test.sv"
	`include "full_76800_5_none_2_test.sv"
	`include "full_76800_5_odd_1_test.sv"
	`include "full_76800_5_odd_2_test.sv"
	`include "full_76800_5_even_1_test.sv"
	`include "full_76800_5_even_2_test.sv"

	`include "full_76800_6_none_1_test.sv"
	`include "full_76800_6_none_2_test.sv"
	`include "full_76800_6_odd_1_test.sv"
	`include "full_76800_6_odd_2_test.sv"
	`include "full_76800_6_even_1_test.sv"
	`include "full_76800_6_even_2_test.sv"

	`include "full_76800_7_none_1_test.sv"
	`include "full_76800_7_none_2_test.sv"
	`include "full_76800_7_odd_1_test.sv"
	`include "full_76800_7_odd_2_test.sv"
	`include "full_76800_7_even_1_test.sv"
	`include "full_76800_7_even_2_test.sv"

	`include "full_76800_8_none_1_test.sv"
	`include "full_76800_8_none_2_test.sv"
	`include "full_76800_8_odd_1_test.sv"
	`include "full_76800_8_odd_2_test.sv"
	`include "full_76800_8_even_1_test.sv"
	`include "full_76800_8_even_2_test.sv"

	`include "full_115200_5_none_1_test.sv"
	`include "full_115200_5_none_2_test.sv"
	`include "full_115200_5_odd_1_test.sv"
	`include "full_115200_5_odd_2_test.sv"
	`include "full_115200_5_even_1_test.sv"
	`include "full_115200_5_even_2_test.sv"

	`include "full_115200_6_none_1_test.sv"
	`include "full_115200_6_none_2_test.sv"
	`include "full_115200_6_odd_1_test.sv"
	`include "full_115200_6_odd_2_test.sv"
	`include "full_115200_6_even_1_test.sv"
	`include "full_115200_6_even_2_test.sv"

	`include "full_115200_7_none_1_test.sv"
	`include "full_115200_7_none_2_test.sv"
	`include "full_115200_7_odd_1_test.sv"
	`include "full_115200_7_odd_2_test.sv"
	`include "full_115200_7_even_1_test.sv"
	`include "full_115200_7_even_2_test.sv"

	`include "full_115200_8_none_1_test.sv"
	`include "full_115200_8_none_2_test.sv"
	`include "full_115200_8_odd_1_test.sv"
	`include "full_115200_8_odd_2_test.sv"
	`include "full_115200_8_even_1_test.sv"
	`include "full_115200_8_even_2_test.sv"

	`include "full_custom_5_none_1_test.sv"
	`include "full_custom_5_none_2_test.sv"
	`include "full_custom_5_odd_1_test.sv"
	`include "full_custom_5_odd_2_test.sv"
	`include "full_custom_5_even_1_test.sv"
	`include "full_custom_5_even_2_test.sv"

	`include "full_custom_6_none_1_test.sv"
	`include "full_custom_6_none_2_test.sv"
	`include "full_custom_6_odd_1_test.sv"
	`include "full_custom_6_odd_2_test.sv"
	`include "full_custom_6_even_1_test.sv"
	`include "full_custom_6_even_2_test.sv"

	`include "full_custom_7_none_1_test.sv"
	`include "full_custom_7_none_2_test.sv"
	`include "full_custom_7_odd_1_test.sv"
	`include "full_custom_7_odd_2_test.sv"
	`include "full_custom_7_even_1_test.sv"
	`include "full_custom_7_even_2_test.sv"

	`include "full_custom_8_none_1_test.sv"
	`include "full_custom_8_none_2_test.sv"
	`include "full_custom_8_odd_1_test.sv"
	`include "full_custom_8_odd_2_test.sv"
	`include "full_custom_8_even_1_test.sv"
	`include "full_custom_8_even_2_test.sv"

	`include "full_dynamic_config_test.sv"
	
	`include "interrupt_parity_error_en_test.sv"
	`include "interrupt_parity_error_dis_test.sv"
	`include "interrupt_rx_empty_en_test.sv"
	`include "interrupt_rx_empty_dis_test.sv"
	`include "interrupt_tx_empty_en_test.sv"
	`include "interrupt_tx_empty_dis_test.sv"
	`include "interrupt_rx_full_en_test.sv"
	`include "interrupt_rx_full_dis_test.sv"
	`include "interrupt_tx_full_en_test.sv"
	`include "interrupt_tx_full_dis_test.sv"

	`include "mismatch_parity_test.sv"
	`include "mismatch_baudrate_test.sv"	
	`include "mismatch_data_width_test.sv"
	`include "mismatch_stop_width_test.sv"

	`include "wr_when_tx_full_test.sv"
endpackage
`endif
